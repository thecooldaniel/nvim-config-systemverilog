package packageExample;

    function void exampleFunc();
        $display("exampleFunc called");
    endfunction

endpackage

