package packageExample;

    function void exampleFunc();
        // Function implementation
        $display("exampleFunc called");
    endfunction

endpackage

